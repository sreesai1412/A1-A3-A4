module demux_32to1 (input [a
