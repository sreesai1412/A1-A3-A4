`include "../lib/mux_16to1.v"

module test;

  reg  [3:0] s;
  reg  i15, i14, i13, i12, i11, i10, i9, i8, i7, i6, i5, i4, i3, i2, i1, i0;
  wire z;

  mux_16to1 mux(
    .s  (s ),
    .i15(i15),   
    .i14(i14),
    .i13(i13),
    .i12(i12),
    .i11(i11),
    .i10(i10),
    .i9 (i9 ),
    .i8 (i8 ),
    .i7 (i7 ),
    .i6 (i6 ),
    .i5 (i5 ),
    .i4 (i4 ),
    .i3 (i3 ),
    .i2 (i2 ),
    .i1 (i1 ),
    .i0 (i0 ),
    .z  (z ));
  
  initial begin
    $monitor($time, ":  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b  %b | %b  %b  %b  %b | %b",
                      i15, i14, i13, i12,i11,i10,i9, i8,i7, i6, i5, i4, i3, i2, i1, i0,s[3], s[2],s[1],s[0],z);
        
    #5 i15  = 0; i14  = 0; i13  = 0; i12  = 0; i11 = 0; i10 = 0; i9 = 0; i8 = 0;  
       i7   = 0; i6   = 0; i5   = 0; i4   = 0; i3  = 0; i2  = 0; i1 = 0; i0 = 0; 
       s[3] = 0; s[2] = 0; s[1] = 0; s[0] = 0;

    #5 i4 = 1; i5 = 1; i2 = 1; s[1] = 1; // 010 select i2
    #5 s[0] = 1; // 0011 select i3
    #5 s[2] = 1; // 0111 select i7
    #5 i7 = 0;
    #5 s[1] = 0; // 0101 select i5
    #5 i15  = 1; s[1] = 1; s[3] = 1; //1111 select i15
    #5 i10 = 1; s[0] = 0; s[2] = 0; // 1010 select i10
  end

// 0000 0
// 0001 1
// 0010 2
// 0011 3
// 0100 4
// 0101 5
// 0110 6
// 0111 7
// 1000 8
// 1001 9
// 1010 10
// 1011 11
// 1100 12
// 1101 13
// 1110 14
// 1111 15
 
endmodule
