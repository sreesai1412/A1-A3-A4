`include "../lib/mux_32to1.v"

module mux32bits_32to1 (
  input  [4:0 ] s,
  input  [31:0] i31, i30, i29, i28, i27, i26, i25, i24, i23,i22, i21, i20, i19, i18, i17, i16,
  input  [31:0] i15, i14, i13, i12, i11, i10, i9, i8, i7,i6, i5, i4, i3, i2, i1, i0,
  output [31:0] z);

mux_32to1 mux0 (.z(z[0 ]), .i31(i31[0 ]), .i30(i30[0 ]), .i29(i29[0 ]), .i28(i28[0 ]), .i27(i27[0 ]), .i26(i26[0 ]), .i25(i25[0 ]), .i24(i24[0 ]), .i23(i23[0 ]), .i22(i22[0 ]), .i21(i21[0 ]), .i20(i20[0 ]), .i19(i19[0 ]), .i18(i18[0 ]), .i17(i17[0 ]), .i16(i16[0 ]), .i15(i15[0 ]), .i14(i14[0 ]), .i13(i13[0 ]), .i12(i12[0 ]), .i11(i11[0 ]), .i10(i10[0 ]), .i9(i9[0 ]), .i8(i8[0 ]), .i7(i7[0 ]), .i6(i6[0 ]), .i5(i5[0 ]), .i4(i4[0 ]), .i3(i3[0 ]), .i2(i2[0 ]), .i1(i1[0 ]), .i0(i0[0 ]), .s(s));

mux_32to1 mux1 (.z(z[1 ]), .i31(i31[1 ]), .i30(i30[1 ]), .i29(i29[1 ]), .i28(i28[1 ]), .i27(i27[1 ]), .i26(i26[1 ]), .i25(i25[1 ]), .i24(i24[1 ]), .i23(i23[1 ]), .i22(i22[1 ]), .i21(i21[1 ]), .i20(i20[1 ]), .i19(i19[1 ]), .i18(i18[1 ]), .i17(i17[1 ]), .i16(i16[1 ]), .i15(i15[1 ]), .i14(i14[1 ]), .i13(i13[1 ]), .i12(i12[1 ]), .i11(i11[1 ]), .i10(i10[1 ]), .i9(i9[1 ]), .i8(i8[1 ]), .i7(i7[1 ]), .i6(i6[1 ]), .i5(i5[1 ]), .i4(i4[1 ]), .i3(i3[1 ]), .i2(i2[1 ]), .i1(i1[1 ]), .i0(i0[1 ]), .s(s));

mux_32to1 mux2 (.z(z[2 ]), .i31(i31[2 ]), .i30(i30[2 ]), .i29(i29[2 ]), .i28(i28[2 ]), .i27(i27[2 ]), .i26(i26[2 ]), .i25(i25[2 ]), .i24(i24[2 ]), .i23(i23[2 ]), .i22(i22[2 ]), .i21(i21[2 ]), .i20(i20[2 ]), .i19(i19[2 ]), .i18(i18[2 ]), .i17(i17[2 ]), .i16(i16[2 ]), .i15(i15[2 ]), .i14(i14[2 ]), .i13(i13[2 ]), .i12(i12[2 ]), .i11(i11[2 ]), .i10(i10[2 ]), .i9(i9[2 ]), .i8(i8[2 ]), .i7(i7[2 ]), .i6(i6[2 ]), .i5(i5[2 ]), .i4(i4[2 ]), .i3(i3[2 ]), .i2(i2[2 ]), .i1(i1[2 ]), .i0(i0[2 ]), .s(s));

mux_32to1 mux3 (.z(z[3 ]), .i31(i31[3 ]), .i30(i30[3 ]), .i29(i29[3 ]), .i28(i28[3 ]), .i27(i27[3 ]), .i26(i26[3 ]), .i25(i25[3 ]), .i24(i24[3 ]), .i23(i23[3 ]), .i22(i22[3 ]), .i21(i21[3 ]), .i20(i20[3 ]), .i19(i19[3 ]), .i18(i18[3 ]), .i17(i17[3 ]), .i16(i16[3 ]), .i15(i15[3 ]), .i14(i14[3 ]), .i13(i13[3 ]), .i12(i12[3 ]), .i11(i11[3 ]), .i10(i10[3 ]), .i9(i9[3 ]), .i8(i8[3 ]), .i7(i7[3 ]), .i6(i6[3 ]), .i5(i5[3 ]), .i4(i4[3 ]), .i3(i3[3 ]), .i2(i2[3 ]), .i1(i1[3 ]), .i0(i0[3 ]), .s(s));

mux_32to1 mux4 (.z(z[4 ]), .i31(i31[4 ]), .i30(i30[4 ]), .i29(i29[4 ]), .i28(i28[4 ]), .i27(i27[4 ]), .i26(i26[4 ]), .i25(i25[4 ]), .i24(i24[4 ]), .i23(i23[4 ]), .i22(i22[4 ]), .i21(i21[4 ]), .i20(i20[4 ]), .i19(i19[4 ]), .i18(i18[4 ]), .i17(i17[4 ]), .i16(i16[4 ]), .i15(i15[4 ]), .i14(i14[4 ]), .i13(i13[4 ]), .i12(i12[4 ]), .i11(i11[4 ]), .i10(i10[4 ]), .i9(i9[4 ]), .i8(i8[4 ]), .i7(i7[4 ]), .i6(i6[4 ]), .i5(i5[4 ]), .i4(i4[4 ]), .i3(i3[4 ]), .i2(i2[4 ]), .i1(i1[4 ]), .i0(i0[4 ]), .s(s));

mux_32to1 mux5 (.z(z[5 ]), .i31(i31[5 ]), .i30(i30[5 ]), .i29(i29[5 ]), .i28(i28[5 ]), .i27(i27[5 ]), .i26(i26[5 ]), .i25(i25[5 ]), .i24(i24[5 ]), .i23(i23[5 ]), .i22(i22[5 ]), .i21(i21[5 ]), .i20(i20[5 ]), .i19(i19[5 ]), .i18(i18[5 ]), .i17(i17[5 ]), .i16(i16[5 ]), .i15(i15[5 ]), .i14(i14[5 ]), .i13(i13[5 ]), .i12(i12[5 ]), .i11(i11[5 ]), .i10(i10[5 ]), .i9(i9[5 ]), .i8(i8[5 ]), .i7(i7[5 ]), .i6(i6[5 ]), .i5(i5[5 ]), .i4(i4[5 ]), .i3(i3[5 ]), .i2(i2[5 ]), .i1(i1[5 ]), .i0(i0[5 ]), .s(s));

mux_32to1 mux6 (.z(z[6 ]), .i31(i31[6 ]), .i30(i30[6 ]), .i29(i29[6 ]), .i28(i28[6 ]), .i27(i27[6 ]), .i26(i26[6 ]), .i25(i25[6 ]), .i24(i24[6 ]), .i23(i23[6 ]), .i22(i22[6 ]), .i21(i21[6 ]), .i20(i20[6 ]), .i19(i19[6 ]), .i18(i18[6 ]), .i17(i17[6 ]), .i16(i16[6 ]), .i15(i15[6 ]), .i14(i14[6 ]), .i13(i13[6 ]), .i12(i12[6 ]), .i11(i11[6 ]), .i10(i10[6 ]), .i9(i9[6 ]), .i8(i8[6 ]), .i7(i7[6 ]), .i6(i6[6 ]), .i5(i5[6 ]), .i4(i4[6 ]), .i3(i3[6 ]), .i2(i2[6 ]), .i1(i1[6 ]), .i0(i0[6 ]), .s(s));

mux_32to1 mux7 (.z(z[7 ]), .i31(i31[7 ]), .i30(i30[7 ]), .i29(i29[7 ]), .i28(i28[7 ]), .i27(i27[7 ]), .i26(i26[7 ]), .i25(i25[7 ]), .i24(i24[7 ]), .i23(i23[7 ]), .i22(i22[7 ]), .i21(i21[7 ]), .i20(i20[7 ]), .i19(i19[7 ]), .i18(i18[7 ]), .i17(i17[7 ]), .i16(i16[7 ]), .i15(i15[7 ]), .i14(i14[7 ]), .i13(i13[7 ]), .i12(i12[7 ]), .i11(i11[7 ]), .i10(i10[7 ]), .i9(i9[7 ]), .i8(i8[7 ]), .i7(i7[7 ]), .i6(i6[7 ]), .i5(i5[7 ]), .i4(i4[7 ]), .i3(i3[7 ]), .i2(i2[7 ]), .i1(i1[7 ]), .i0(i0[7 ]), .s(s));

mux_32to1 mux8 (.z(z[8 ]), .i31(i31[8 ]), .i30(i30[8 ]), .i29(i29[8 ]), .i28(i28[8 ]), .i27(i27[8 ]), .i26(i26[8 ]), .i25(i25[8 ]), .i24(i24[8 ]), .i23(i23[8 ]), .i22(i22[8 ]), .i21(i21[8 ]), .i20(i20[8 ]), .i19(i19[8 ]), .i18(i18[8 ]), .i17(i17[8 ]), .i16(i16[8 ]), .i15(i15[8 ]), .i14(i14[8 ]), .i13(i13[8 ]), .i12(i12[8 ]), .i11(i11[8 ]), .i10(i10[8 ]), .i9(i9[8 ]), .i8(i8[8 ]), .i7(i7[8 ]), .i6(i6[8 ]), .i5(i5[8 ]), .i4(i4[8 ]), .i3(i3[8 ]), .i2(i2[8 ]), .i1(i1[8 ]), .i0(i0[8 ]), .s(s));

mux_32to1 mux9 (.z(z[9 ]), .i31(i31[9 ]), .i30(i30[9 ]), .i29(i29[9 ]), .i28(i28[9 ]), .i27(i27[9 ]), .i26(i26[9 ]), .i25(i25[9 ]), .i24(i24[9 ]), .i23(i23[9 ]), .i22(i22[9 ]), .i21(i21[9 ]), .i20(i20[9 ]), .i19(i19[9 ]), .i18(i18[9 ]), .i17(i17[9 ]), .i16(i16[9 ]), .i15(i15[9 ]), .i14(i14[9 ]), .i13(i13[9 ]), .i12(i12[9 ]), .i11(i11[9 ]), .i10(i10[9 ]), .i9(i9[9 ]), .i8(i8[9 ]), .i7(i7[9 ]), .i6(i6[9 ]), .i5(i5[9 ]), .i4(i4[9 ]), .i3(i3[9 ]), .i2(i2[9 ]), .i1(i1[9 ]), .i0(i0[9 ]), .s(s));

mux_32to1 mux10(.z(z[10]), .i31(i31[10]), .i30(i30[10]), .i29(i29[10]), .i28(i28[10]), .i27(i27[10]), .i26(i26[10]), .i25(i25[10]), .i24(i24[10]), .i23(i23[10]), .i22(i22[10]), .i21(i21[10]), .i20(i20[10]), .i19(i19[10]), .i18(i18[10]), .i17(i17[10]), .i16(i16[10]), .i15(i15[10]), .i14(i14[10]), .i13(i13[10]), .i12(i12[10]), .i11(i11[10]), .i10(i10[10]), .i9(i9[10]), .i8(i8[10]), .i7(i7[10]), .i6(i6[10]), .i5(i5[10]), .i4(i4[10]), .i3(i3[10]), .i2(i2[10]), .i1(i1[10]), .i0(i0[10]), .s(s));

mux_32to1 mux11(.z(z[11]), .i31(i31[11]), .i30(i30[11]), .i29(i29[11]), .i28(i28[11]), .i27(i27[11]), .i26(i26[11]), .i25(i25[11]), .i24(i24[11]), .i23(i23[11]), .i22(i22[11]), .i21(i21[11]), .i20(i20[11]), .i19(i19[11]), .i18(i18[11]), .i17(i17[11]), .i16(i16[11]), .i15(i15[11]), .i14(i14[11]), .i13(i13[11]), .i12(i12[11]), .i11(i11[11]), .i10(i10[11]), .i9(i9[11]), .i8(i8[11]), .i7(i7[11]), .i6(i6[11]), .i5(i5[11]), .i4(i4[11]), .i3(i3[11]), .i2(i2[11]), .i1(i1[11]), .i0(i0[11]), .s(s));

mux_32to1 mux12(.z(z[12]), .i31(i31[12]), .i30(i30[12]), .i29(i29[12]), .i28(i28[12]), .i27(i27[12]), .i26(i26[12]), .i25(i25[12]), .i24(i24[12]), .i23(i23[12]), .i22(i22[12]), .i21(i21[12]), .i20(i20[12]), .i19(i19[12]), .i18(i18[12]), .i17(i17[12]), .i16(i16[12]), .i15(i15[12]), .i14(i14[12]), .i13(i13[12]), .i12(i12[12]), .i11(i11[12]), .i10(i10[12]), .i9(i9[12]), .i8(i8[12]), .i7(i7[12]), .i6(i6[12]), .i5(i5[12]), .i4(i4[12]), .i3(i3[12]), .i2(i2[12]), .i1(i1[12]), .i0(i0[12]), .s(s));

mux_32to1 mux13(.z(z[13]), .i31(i31[13]), .i30(i30[13]), .i29(i29[13]), .i28(i28[13]), .i27(i27[13]), .i26(i26[13]), .i25(i25[13]), .i24(i24[13]), .i23(i23[13]), .i22(i22[13]), .i21(i21[13]), .i20(i20[13]), .i19(i19[13]), .i18(i18[13]), .i17(i17[13]), .i16(i16[13]), .i15(i15[13]), .i14(i14[13]), .i13(i13[13]), .i12(i12[13]), .i11(i11[13]), .i10(i10[13]), .i9(i9[13]), .i8(i8[13]), .i7(i7[13]), .i6(i6[13]), .i5(i5[13]), .i4(i4[13]), .i3(i3[13]), .i2(i2[13]), .i1(i1[13]), .i0(i0[13]), .s(s));

mux_32to1 mux14(.z(z[14]), .i31(i31[14]), .i30(i30[14]), .i29(i29[14]), .i28(i28[14]), .i27(i27[14]), .i26(i26[14]), .i25(i25[14]), .i24(i24[14]), .i23(i23[14]), .i22(i22[14]), .i21(i21[14]), .i20(i20[14]), .i19(i19[14]), .i18(i18[14]), .i17(i17[14]), .i16(i16[14]), .i15(i15[14]), .i14(i14[14]), .i13(i13[14]), .i12(i12[14]), .i11(i11[14]), .i10(i10[14]), .i9(i9[14]), .i8(i8[14]), .i7(i7[14]), .i6(i6[14]), .i5(i5[14]), .i4(i4[14]), .i3(i3[14]), .i2(i2[14]), .i1(i1[14]), .i0(i0[14]), .s(s));

mux_32to1 mux15(.z(z[15]), .i31(i31[15]), .i30(i30[15]), .i29(i29[15]), .i28(i28[15]), .i27(i27[15]), .i26(i26[15]), .i25(i25[15]), .i24(i24[15]), .i23(i23[15]), .i22(i22[15]), .i21(i21[15]), .i20(i20[15]), .i19(i19[15]), .i18(i18[15]), .i17(i17[15]), .i16(i16[15]), .i15(i15[15]), .i14(i14[15]), .i13(i13[15]), .i12(i12[15]), .i11(i11[15]), .i10(i10[15]), .i9(i9[15]), .i8(i8[15]), .i7(i7[15]), .i6(i6[15]), .i5(i5[15]), .i4(i4[15]), .i3(i3[15]), .i2(i2[15]), .i1(i1[15]), .i0(i0[15]), .s(s));

mux_32to1 mux16(.z(z[16]), .i31(i31[16]), .i30(i30[16]), .i29(i29[16]), .i28(i28[16]), .i27(i27[16]), .i26(i26[16]), .i25(i25[16]), .i24(i24[16]), .i23(i23[16]), .i22(i22[16]), .i21(i21[16]), .i20(i20[16]), .i19(i19[16]), .i18(i18[16]), .i17(i17[16]), .i16(i16[16]), .i15(i15[16]), .i14(i14[16]), .i13(i13[16]), .i12(i12[16]), .i11(i11[16]), .i10(i10[16]), .i9(i9[16]), .i8(i8[16]), .i7(i7[16]), .i6(i6[16]), .i5(i5[16]), .i4(i4[16]), .i3(i3[16]), .i2(i2[16]), .i1(i1[16]), .i0(i0[16]), .s(s));

mux_32to1 mux17(.z(z[17]), .i31(i31[17]), .i30(i30[17]), .i29(i29[17]), .i28(i28[17]), .i27(i27[17]), .i26(i26[17]), .i25(i25[17]), .i24(i24[17]), .i23(i23[17]), .i22(i22[17]), .i21(i21[17]), .i20(i20[17]), .i19(i19[17]), .i18(i18[17]), .i17(i17[17]), .i16(i16[17]), .i15(i15[17]), .i14(i14[17]), .i13(i13[17]), .i12(i12[17]), .i11(i11[17]), .i10(i10[17]), .i9(i9[17]), .i8(i8[17]), .i7(i7[17]), .i6(i6[17]), .i5(i5[17]), .i4(i4[17]), .i3(i3[17]), .i2(i2[17]), .i1(i1[17]), .i0(i0[17]), .s(s));

mux_32to1 mux18(.z(z[18]), .i31(i31[18]), .i30(i30[18]), .i29(i29[18]), .i28(i28[18]), .i27(i27[18]), .i26(i26[18]), .i25(i25[18]), .i24(i24[18]), .i23(i23[18]), .i22(i22[18]), .i21(i21[18]), .i20(i20[18]), .i19(i19[18]), .i18(i18[18]), .i17(i17[18]), .i16(i16[18]), .i15(i15[18]), .i14(i14[18]), .i13(i13[18]), .i12(i12[18]), .i11(i11[18]), .i10(i10[18]), .i9(i9[18]), .i8(i8[18]), .i7(i7[18]), .i6(i6[18]), .i5(i5[18]), .i4(i4[18]), .i3(i3[18]), .i2(i2[18]), .i1(i1[18]), .i0(i0[18]), .s(s));

mux_32to1 mux19(.z(z[19]), .i31(i31[19]), .i30(i30[19]), .i29(i29[19]), .i28(i28[19]), .i27(i27[19]), .i26(i26[19]), .i25(i25[19]), .i24(i24[19]), .i23(i23[19]), .i22(i22[19]), .i21(i21[19]), .i20(i20[19]), .i19(i19[19]), .i18(i18[19]), .i17(i17[19]), .i16(i16[19]), .i15(i15[19]), .i14(i14[19]), .i13(i13[19]), .i12(i12[19]), .i11(i11[19]), .i10(i10[19]), .i9(i9[19]), .i8(i8[19]), .i7(i7[19]), .i6(i6[19]), .i5(i5[19]), .i4(i4[19]), .i3(i3[19]), .i2(i2[19]), .i1(i1[19]), .i0(i0[19]), .s(s));

mux_32to1 mux20(.z(z[20]), .i31(i31[20]), .i30(i30[20]), .i29(i29[20]), .i28(i28[20]), .i27(i27[20]), .i26(i26[20]), .i25(i25[20]), .i24(i24[20]), .i23(i23[20]), .i22(i22[20]), .i21(i21[20]), .i20(i20[20]), .i19(i19[20]), .i18(i18[20]), .i17(i17[20]), .i16(i16[20]), .i15(i15[20]), .i14(i14[20]), .i13(i13[20]), .i12(i12[20]), .i11(i11[20]), .i10(i10[20]), .i9(i9[20]), .i8(i8[20]), .i7(i7[20]), .i6(i6[20]), .i5(i5[20]), .i4(i4[20]), .i3(i3[20]), .i2(i2[20]), .i1(i1[20]), .i0(i0[20]), .s(s));

mux_32to1 mux21(.z(z[21]), .i31(i31[21]), .i30(i30[21]), .i29(i29[21]), .i28(i28[21]), .i27(i27[21]), .i26(i26[21]), .i25(i25[21]), .i24(i24[21]), .i23(i23[21]), .i22(i22[21]), .i21(i21[21]), .i20(i20[21]), .i19(i19[21]), .i18(i18[21]), .i17(i17[21]), .i16(i16[21]), .i15(i15[21]), .i14(i14[21]), .i13(i13[21]), .i12(i12[21]), .i11(i11[21]), .i10(i10[21]), .i9(i9[21]), .i8(i8[21]), .i7(i7[21]), .i6(i6[21]), .i5(i5[21]), .i4(i4[21]), .i3(i3[21]), .i2(i2[21]), .i1(i1[21]), .i0(i0[21]), .s(s));

mux_32to1 mux22(.z(z[22]), .i31(i31[22]), .i30(i30[22]), .i29(i29[22]), .i28(i28[22]), .i27(i27[22]), .i26(i26[22]), .i25(i25[22]), .i24(i24[22]), .i23(i23[22]), .i22(i22[22]), .i21(i21[22]), .i20(i20[22]), .i19(i19[22]), .i18(i18[22]), .i17(i17[22]), .i16(i16[22]), .i15(i15[22]), .i14(i14[22]), .i13(i13[22]), .i12(i12[22]), .i11(i11[22]), .i10(i10[22]), .i9(i9[22]), .i8(i8[22]), .i7(i7[22]), .i6(i6[22]), .i5(i5[22]), .i4(i4[22]), .i3(i3[22]), .i2(i2[22]), .i1(i1[22]), .i0(i0[22]), .s(s));


mux_32to1 mux23(.z(z[23]), .i31(i31[23]), .i30(i30[23]), .i29(i29[23]), .i28(i28[23]), .i27(i27[23]), .i26(i26[23]), .i25(i25[23]), .i24(i24[23]), .i23(i23[23]), .i22(i22[23]), .i21(i21[23]), .i20(i20[23]), .i19(i19[23]), .i18(i18[23]), .i17(i17[23]), .i16(i16[23]), .i15(i15[23]), .i14(i14[23]), .i13(i13[23]), .i12(i12[23]), .i11(i11[23]), .i10(i10[23]), .i9(i9[23]), .i8(i8[23]), .i7(i7[23]), .i6(i6[23]), .i5(i5[23]), .i4(i4[23]), .i3(i3[23]), .i2(i2[23]), .i1(i1[23]), .i0(i0[23]), .s(s));

mux_32to1 mux24(.z(z[24]), .i31(i31[24]), .i30(i30[24]), .i29(i29[24]), .i28(i28[24]), .i27(i27[24]), .i26(i26[24]), .i25(i25[24]), .i24(i24[24]), .i23(i23[24]), .i22(i22[24]), .i21(i21[24]), .i20(i20[24]), .i19(i19[24]), .i18(i18[24]), .i17(i17[24]), .i16(i16[24]), .i15(i15[24]), .i14(i14[24]), .i13(i13[24]), .i12(i12[24]), .i11(i11[24]), .i10(i10[24]), .i9(i9[24]), .i8(i8[24]), .i7(i7[24]), .i6(i6[24]), .i5(i5[24]), .i4(i4[24]), .i3(i3[24]), .i2(i2[24]), .i1(i1[24]), .i0(i0[24]), .s(s));

mux_32to1 mux25(.z(z[25]), .i31(i31[25]), .i30(i30[25]), .i29(i29[25]), .i28(i28[25]), .i27(i27[25]), .i26(i26[25]), .i25(i25[25]), .i24(i24[25]), .i23(i23[25]), .i22(i22[25]), .i21(i21[25]), .i20(i20[25]), .i19(i19[25]), .i18(i18[25]), .i17(i17[25]), .i16(i16[25]), .i15(i15[25]), .i14(i14[25]), .i13(i13[25]), .i12(i12[25]), .i11(i11[25]), .i10(i10[25]), .i9(i9[25]), .i8(i8[25]), .i7(i7[25]), .i6(i6[25]), .i5(i5[25]), .i4(i4[25]), .i3(i3[25]), .i2(i2[25]), .i1(i1[25]), .i0(i0[25]), .s(s));

mux_32to1 mux26(.z(z[26]), .i31(i31[26]), .i30(i30[26]), .i29(i29[26]), .i28(i28[26]), .i27(i27[26]), .i26(i26[26]), .i25(i25[26]), .i24(i24[26]), .i23(i23[26]), .i22(i22[26]), .i21(i21[26]), .i20(i20[26]), .i19(i19[26]), .i18(i18[26]), .i17(i17[26]), .i16(i16[26]), .i15(i15[26]), .i14(i14[26]), .i13(i13[26]), .i12(i12[26]), .i11(i11[26]), .i10(i10[26]), .i9(i9[26]), .i8(i8[26]), .i7(i7[26]), .i6(i6[26]), .i5(i5[26]), .i4(i4[26]), .i3(i3[26]), .i2(i2[26]), .i1(i1[26]), .i0(i0[26]), .s(s));

mux_32to1 mux27(.z(z[27]), .i31(i31[27]), .i30(i30[27]), .i29(i29[27]), .i28(i28[27]), .i27(i27[27]), .i26(i26[27]), .i25(i25[27]), .i24(i24[27]), .i23(i23[27]), .i22(i22[27]), .i21(i21[27]), .i20(i20[27]), .i19(i19[27]), .i18(i18[27]), .i17(i17[27]), .i16(i16[27]), .i15(i15[27]), .i14(i14[27]), .i13(i13[27]), .i12(i12[27]), .i11(i11[27]), .i10(i10[27]), .i9(i9[27]), .i8(i8[27]), .i7(i7[27]), .i6(i6[27]), .i5(i5[27]), .i4(i4[27]), .i3(i3[27]), .i2(i2[27]), .i1(i1[27]), .i0(i0[27]), .s(s));

mux_32to1 mux28(.z(z[28]), .i31(i31[28]), .i30(i30[28]), .i29(i29[28]), .i28(i28[28]), .i27(i27[28]), .i26(i26[28]), .i25(i25[28]), .i24(i24[28]), .i23(i23[28]), .i22(i22[28]), .i21(i21[28]), .i20(i20[28]), .i19(i19[28]), .i18(i18[28]), .i17(i17[28]), .i16(i16[28]), .i15(i15[28]), .i14(i14[28]), .i13(i13[28]), .i12(i12[28]), .i11(i11[28]), .i10(i10[28]), .i9(i9[28]), .i8(i8[28]), .i7(i7[28]), .i6(i6[28]), .i5(i5[28]), .i4(i4[28]), .i3(i3[28]), .i2(i2[28]), .i1(i1[28]), .i0(i0[28]), .s(s));

mux_32to1 mux29(.z(z[29]), .i31(i31[29]), .i30(i30[29]), .i29(i29[29]), .i28(i28[29]), .i27(i27[29]), .i26(i26[29]), .i25(i25[29]), .i24(i24[29]), .i23(i23[29]), .i22(i22[29]), .i21(i21[29]), .i20(i20[29]), .i19(i19[29]), .i18(i18[29]), .i17(i17[29]), .i16(i16[29]), .i15(i15[29]), .i14(i14[29]), .i13(i13[29]), .i12(i12[29]), .i11(i11[29]), .i10(i10[29]), .i9(i9[29]), .i8(i8[29]), .i7(i7[29]), .i6(i6[29]), .i5(i5[29]), .i4(i4[29]), .i3(i3[29]), .i2(i2[29]), .i1(i1[29]), .i0(i0[29]), .s(s));

mux_32to1 mux30(.z(z[30]), .i31(i31[30]), .i30(i30[30]), .i29(i29[30]), .i28(i28[30]), .i27(i27[30]), .i26(i26[30]), .i25(i25[30]), .i24(i24[30]), .i23(i23[30]), .i22(i22[30]), .i21(i21[30]), .i20(i20[30]), .i19(i19[30]), .i18(i18[30]), .i17(i17[30]), .i16(i16[30]), .i15(i15[30]), .i14(i14[30]), .i13(i13[30]), .i12(i12[30]), .i11(i11[30]), .i10(i10[30]), .i9(i9[30]), .i8(i8[30]), .i7(i7[30]), .i6(i6[30]), .i5(i5[30]), .i4(i4[30]), .i3(i3[30]), .i2(i2[30]), .i1(i1[30]), .i0(i0[30]), .s(s));

mux_32to1 mux31(.z(z[31]), .i31(i31[31]), .i30(i30[31]), .i29(i29[31]), .i28(i28[31]), .i27(i27[31]), .i26(i26[31]), .i25(i25[31]), .i24(i24[31]), .i23(i23[31]), .i22(i22[31]), .i21(i21[31]), .i20(i20[31]), .i19(i19[31]), .i18(i18[31]), .i17(i17[31]), .i16(i16[31]), .i15(i15[31]), .i14(i14[31]), .i13(i13[31]), .i12(i12[31]), .i11(i11[31]), .i10(i10[31]), .i9(i9[31]), .i8(i8[31]), .i7(i7[31]), .i6(i6[31]), .i5(i5[31]), .i4(i4[31]), .i3(i3[31]), .i2(i2[31]), .i1(i1[31]), .i0(i0[31]), .s(s));

endmodule
