module alu_control ( 
  input [5:0] funct,
  input [1:0] alu_op,
  output [3:0] aluctrl);

  always @(*) begin
    case(funct
  end

endmodule
